module logicgates(a,b,andgate,orgate,xorgate,nandgate,norgate,xnorgate,notgate);
input a,b;
output andgate,orgate,xorgate,nandgate,norgate,xnorgate,notgate;
and (andgate,a,b);
or (orgate,a,b);
xor (xorgate,a,b);
nand (nandgate,a,b);  
nor (norgate,a,b);
xnor (xnorgate,a,b);
not (notgate,a);
endmodule
